module temp_controle (clk_controle, reset, arm, limp, hab);   
    input clk_controle, reset;
    output bit arm, limp, hab;
endmodule
