module contDec(clk_in, reset, clk_out);
  input clk_in, reset;
  output bit clk_out;
endmodule
