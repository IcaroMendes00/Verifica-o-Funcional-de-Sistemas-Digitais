module cont_BCD (clk_amostra, reset, limp, hab, cont_3, cont_2, cont_1, cont_0  );   
    input clk_amostra, reset, limp, hab;
    output logic [3:0] cont_3, cont_2, cont_1, cont_0;
endmodule
